/////////////////////////////////////////////////////////////////////////
//                                                                     //
//  Modulename  :  IB.sv                                               //
//                                                                     //
//  Description :  Issue Buffer. Buffering the issued instructions to  //
//                 different types of Function Units, and route them   //
//                 to a specific Function Unit based on availibility.  //
//                                                                     //
/////////////////////////////////////////////////////////////////////////

module IB #(
    parameter   C_IS_NUM        =   `IS_NUM     ,
    parameter   C_ALU_BASE      =   `ALU_BASE   , 
    parameter   C_MULT_BASE     =   `MULT_BASE  , 
    parameter   C_BR_BASE       =   `BR_BASE    , 
    parameter   C_LOAD_BASE     =   `LOAD_BASE  , 
    parameter   C_STORE_BASE    =   `STORE_BASE , 
    parameter   C_FU_NUM        =   `FU_NUM     
) (
    input   logic                       clk_i           ,   //  Clock
    input   logic                       rst_i           ,   //  Reset
    output  IB_RS                       ib_rs_o         ,
    input   RS_IB   [C_IS_NUM-1:0]      rs_ib_i         ,
    output  IB_FU   [C_FU_NUM-1:0]      ib_fu_o         
);

// ====================================================================
// Local Parameters Declarations Start
// ====================================================================

// ====================================================================
// Local Parameters Declarations End
// ====================================================================

// ====================================================================
// Signal Declarations Start
// ====================================================================

// ====================================================================
// Signal Declarations End
// ====================================================================

// ====================================================================
// Module Instantiations Start
// ====================================================================
// --------------------------------------------------------------------
// Module name  :   sub_module_name
// Description  :   sub module function
// --------------------------------------------------------------------


// --------------------------------------------------------------------


// ====================================================================
// Module Instantiations End
// ====================================================================

// ====================================================================
// RTL Logic Start
// ====================================================================

// --------------------------------------------------------------------
// Logic Divider
// --------------------------------------------------------------------

// ====================================================================
// RTL Logic End
// ====================================================================


endmodule
