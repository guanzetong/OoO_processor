
module AMT #(
    parameter C_RT_NUM            = `RT_NUM,
    parameter C_MT_ENTRY = `MT_ENTRY,
    parameter C_TAG_IDX_WIDTH = `TAG_IDX_WIDTH
)(
    input   logic           clk_i,
    input   logic           rst_i,
    input   logic                                   rollback_i, 
    input   DP_AMT   [C_RT_NUM-1:0]      dp_amt_i, 
   
    output  AMT_OUTPUT   [C_MT_ENTRY-1:0] amt_o

);

    AMT_ENTRY  [C_RT_NUM- 1:0] amt_entry;

    always_comb begin
        if (rollback_i) begin
            for (int i=0; i<C_MT_ENTRY; i++) begin
                if (dp_amt_i[0].wr_en && dp_amt_i[0].rd == i) begin
                    amt_o[i].amt_tag = dp_amt_i[0].tag_old;
                end else if (dp_amt_i[1].wr_en && dp_amt_i[1].rd == i) begin
                    amt_o[i].amt_tag = dp_amt_i[1].tag_old;
                end else begin
                    amt_o[i].amt_tag = amt_entry[i].amt_tag;
                end
            end
        end else begin
            for (int i=0; i<C_MT_ENTRY; i++) begin
                amt_o[i].amt_tag = amt_entry[i].amt_tag;
            end
        end
            
    end

    always_ff @(posedge clk_i) begin
        if (rst_i) begin
            for(int i=0; i<C_MT_ENTRY; i++) begin
                amt_entry[i].amt_tag <= i;
            end
        end else begin
            for (int i=0; i<C_MT_ENTRY; i++) begin
                for (int j=0; j<C_RT_NUM; j++) begin
                    if (dp_amt_i[j].wr_en && dp_amt_i[j].rd == i) begin
                        amt_entry[dp_amt_i[j].rd].amt_tag <= dp_amt_i[j].tag_old;
                    end else begin
                    end
                end
            end
        end
    end
    
endmodule