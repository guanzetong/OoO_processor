/////////////////////////////////////////////////////////////////////////
//                                                                     //
//  Modulename  :  template.sv                                         //
//                                                                     //
//  Description :  template                                            // 
//                                                                     //
/////////////////////////////////////////////////////////////////////////

module module_name #(
    parameter   C_PARAM     =   0                   //  A place holder. Delete it.
) (
    input   logic               clk_i           ,   //  Clock
    input   logic               rst_i           ,   //  Reset
    output  logic               dummy               //  A place holder. Delete it.
);

// ====================================================================
// Local Parameters Declarations Start
// ====================================================================

// ====================================================================
// Local Parameters Declarations End
// ====================================================================

// ====================================================================
// Signal Declarations Start
// ====================================================================

// ====================================================================
// Signal Declarations End
// ====================================================================

// ====================================================================
// Module Instantiations Start
// ====================================================================
// --------------------------------------------------------------------
// Module name  :   sub_module_name
// Description  :   sub module function
// --------------------------------------------------------------------


// --------------------------------------------------------------------


// ====================================================================
// Module Instantiations End
// ====================================================================

// ====================================================================
// RTL Logic Start
// ====================================================================

// --------------------------------------------------------------------
// Logic Divider
// --------------------------------------------------------------------

// ====================================================================
// RTL Logic End
// ====================================================================


endmodule
