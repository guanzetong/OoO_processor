/////////////////////////////////////////////////////////////////////////
//                                                                     //
//  Modulename  :  VFL_sim.sv                                          //
//                                                                     //
//  Description :  VFL_sim                                             // 
//                                                                     //
/////////////////////////////////////////////////////////////////////////

module VFL_sim #(
    parameter   C_RT_NUM            =   `RT_NUM         ,
    parameter   C_ARCH_REG_NUM      =   `ARCH_REG_NUM   ,
    parameter   C_PHY_REG_NUM       =   `PHY_REG_NUM    ,
    parameter   C_FL_ENTRY_NUM      =   C_PHY_REG_NUM - C_PHY_REG_NUM
) (
    input   logic                           clk_i       ,   //  Clock
    input   logic                           rst_i       ,   //  Reset
    input   ROB_VFL [C_RT_NUM-1:0]          rob_vfl_i   ,
    output  VFL     [C_FL_ENTRY_NUM-1:0]    vlf_o       ,
    input   logic                           roll_back_i 
);

// ====================================================================
// Local Parameters Declarations Start
// ====================================================================

// ====================================================================
// Local Parameters Declarations End
// ====================================================================

// ====================================================================
// Signal Declarations Start
// ====================================================================

// ====================================================================
// Signal Declarations End
// ====================================================================

// ====================================================================
// Module Instantiations Start
// ====================================================================
// --------------------------------------------------------------------
// Module name  :   sub_module_name
// Description  :   sub module function
// --------------------------------------------------------------------


// --------------------------------------------------------------------


// ====================================================================
// Module Instantiations End
// ====================================================================

// ====================================================================
// RTL Logic Start
// ====================================================================

// --------------------------------------------------------------------
// Logic Divider
// --------------------------------------------------------------------
    task victim_freelist_init();
        begin
            for (int unsigned entry_idx = 0; entry_idx < C_FL_ENTRY_NUM; entry_idx++) begin
                fl_entry.tag    =   entry_idx + C_ARCH_REG_NUM - 1;
                freelist.push_back(fl_entry);
            end
        end
    endtask

    initial begin
        victim_freelist_init();
        victim_freelist_run();
    end
// ====================================================================
// RTL Logic End
// ====================================================================


endmodule
