module test_tb;
    initial begin
        // #50;
        $finish;
    end
    
endmodule