module Freelist_tb (
  ports
);
  
endmodule