/////////////////////////////////////////////////////////////////////////
//                                                                     //
//  Modulename  :  VFL.sv                                              //
//                                                                     //
//  Description :  Victim Freelist                                     // 
//                                                                     //
/////////////////////////////////////////////////////////////////////////

module VFL #(
    parameter   C_RT_NUM    =   `RT_NUM
) (
    input   logic                   clk_i           ,   //  Clock
    input   logic                   rst_i           ,   //  Reset
    input   logic   [C_RT_NUM-1:0]  rob_vfl_i       ,
);

// ====================================================================
// Local Parameters Declarations Start
// ====================================================================

// ====================================================================
// Local Parameters Declarations End
// ====================================================================

// ====================================================================
// Signal Declarations Start
// ====================================================================

// ====================================================================
// Signal Declarations End
// ====================================================================

// ====================================================================
// Module Instantiations Start
// ====================================================================
// --------------------------------------------------------------------
// Module name  :   sub_module_name
// Description  :   sub module function
// --------------------------------------------------------------------


// --------------------------------------------------------------------


// ====================================================================
// Module Instantiations End
// ====================================================================

// ====================================================================
// RTL Logic Start
// ====================================================================

// --------------------------------------------------------------------
// Logic Divider
// --------------------------------------------------------------------

// ====================================================================
// RTL Logic End
// ====================================================================


endmodule
